`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:37:25 03/31/2018 
// Design Name: 
// Module Name:    Switch24To12 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Switch24To12(
	input [3:0] CLH,CLL,
	input CP,nCR,Ctrl
    );
	 //Hour[7:4],Hour[3:0],CP1,nCR,Ctrl24To12
	 
	 always@()


endmodule
